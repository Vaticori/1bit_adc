** sch_path: /headless/Documents/1bit_adc/capacitative_dac.sch
**.subckt capacitative_dac OUT SAR_SEL_1 CLK SAR_SEL_0 SAR_SEL_2 VO_CUR SIN
*.opin OUT
*.ipin SAR_SEL_1
*.ipin CLK
*.ipin SAR_SEL_0
*.ipin SAR_SEL_2
*.opin VO_CUR
*.ipin SIN
XM7 net4 CLK net5 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net6 net7 VSS VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 VREF SAR_SEL_1 S1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=150 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VSS SAR_SEL_0 S0 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=100 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 VSS SAR_SEL_1 S1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=100 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 VSS SAR_SEL_2 S2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=100 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 VREF SAR_SEL_2 S2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=150 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 VREF SAR_SEL_0 S0 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=150 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC3 OUT S2 sky130_fd_pr__cap_mim_m3_1 W=5 L=1 MF=1 m=1
XC5 OUT S2 sky130_fd_pr__cap_mim_m3_1 W=5 L=1 MF=1 m=1
XC6 OUT S2 sky130_fd_pr__cap_mim_m3_1 W=5 L=1 MF=1 m=1
XC7 OUT S1 sky130_fd_pr__cap_mim_m3_1 W=5 L=1 MF=1 m=1
XC8 OUT S1 sky130_fd_pr__cap_mim_m3_1 W=5 L=1 MF=1 m=1
XC9 OUT S0 sky130_fd_pr__cap_mim_m3_1 W=5 L=1 MF=1 m=1
XC10 OUT S2 sky130_fd_pr__cap_mim_m3_1 W=5 L=1 MF=1 m=1
XC11 OUT S2 sky130_fd_pr__cap_mim_m3_1 W=5 L=1 MF=1 m=1
x1 SIN VGND VNB VPB VPWR OUT_BUFF sky130_fd_sc_hd__buf_1
XR1 net8 VDD VSS sky130_fd_pr__res_high_po_0p35 L=0.35 mult=1 m=1
XM9 net9 CURR_ON net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=150 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net8 CURR_ON net10 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=150 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 net3 VSS net1 VSS sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net1 VC_OUT net2 VSS sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net3 net2 VREF VREF sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 VREF net2 net2 VREF sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
VO_CURR net9 VO_CUR 0
.save i(vo_curr)
XC1 VC_OUT VC_IN sky130_fd_pr__cap_mim_m3_1 W=5 L=1 MF=1 m=1
XM15 VC_IN CLK OUT_BUFF VSS sky130_fd_pr__nfet_01v8 L=0.15 W=150 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
VO_CURR1 net10 VSS 0
.save i(vo_curr1)
VO_CURR2 net8 CURR_ON 0
.save i(vo_curr2)
**** begin user architecture code



.option savecurrents

.param vdd=1.8
.param clk=300n
.param settle_time=0.2u
VVDD VDD 0 DC {vdd}
*VCLK CLK 0 PULSE(0 1.8 0 1n 1n 40n 80n)
VVSS VSS 0 DC 0

VVREF VREF 0 DC 1.8

*VSAR_SEL_2 SAR_SEL_2 0  PULSE(0 1.8 0 1n 1n 40n 80n)
*VSAR_SEL_1 SAR_SEL_1 0  PULSE(0 1.8 0 1n 1n 80n 160n)
*VSAR_SEL_0 SAR_SEL_0 0  PULSE(0 1.8 0 1n 1n 160n 320n)

VCLK CLK 0 PULSE(0 1.8 0 1n 1n 20n {settle_time})
VSAR_SEL_2 SAR_SEL_2 0  PULSE(0 1.8 0 1n 1n {2*settle_time} {4*settle_time})
VSAR_SEL_1 SAR_SEL_1 0  PULSE(0 1.8 0 1n 1n {4*settle_time} {8*settle_time})
VSAR_SEL_0 SAR_SEL_0 0  PULSE(0 1.8 0 1n 1n {8*settle_time} {16*settle_time})

VSIN SIN 0 PULSE(0 1.8 0 1n 1n 40n 80n)
VEN EN 0 pwl(0 0  8u 0  8.1u 1.8  16u 1.8  16.1u 0  24u 0  24.1u 1.8  32u 1.8)


.tran 2n 7000n
.control

save all
echo TRAN
run
write 3bit_dac.raw all

.endc
.end



** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include /foss/pdks/sky130A/libs.tech/xschem/sky130_stdcells/

**** end user architecture code
**.ends
.GLOBAL VSS
.GLOBAL VREF
.GLOBAL VDD
.end
