** sch_path: /headless/Documents/1bit_adc/test_three_bit_adc.sch
**.subckt test_three_bit_adc RESET done add sel_wire2,sel_wire1,sel_wire0 CLK
*.ipin RESET
*.opin done
*.ipin add
*.opin sel_wire2,sel_wire1,sel_wire0
*.ipin CLK
ADUT [CLK sel_wire2 sel_wire1 sel_wire0 add RESET done] three_bit_adc
ACOMP [ CLK ] [ clk1 ] adc_buff
A1 [ add ] [ add1 ] adc_buff
ACOMP2 [ RESET ] [ reset1 ] adc_buff
**** begin user architecture code


.param vdd=1.8
VVDD VDD 0 DC {vdd}
VCLK CLK 0 PULSE(0 1.8 0   1n 1n 40n 80n)
Vadd add 0 PULSE(0 1.8 0   1n 1n 10n 80n)
VRESET RESET 0 PULSE(0 1.8 0 1n 1n 40n 800n)
VVSS VSS 0 DC 0
.tran 2n 7000n
.control

save all
echo TRAN
run
write 3bit_adc.raw all
.endc
.end




**** end user architecture code
**.ends

* expanding   symbol:  /headless/Documents/1bit_adc/three_bit_adc.sym # of pins=5
** sym_path: /headless/Documents/1bit_adc/three_bit_adc.sym
** sch_path: /headless/Documents/1bit_adc/three_bit_adc.sch
.subckt three_bit_adc clk sel_wire2 sel_wire1 sel_wire0 add reset done
*.ipin clk
*.ipin reset
*.opin done
*.ipin add
*.opin sel_wire2,sel_wire1,sel_wire0
.ends

**** begin user architecture code
.model three_bit_Adc d_cosim simulation="./three_bit_adc.so"
.model adc_buff adc_bridge in_low=0 in_high=1.1
**** end user architecture code
.end
