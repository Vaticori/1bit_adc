** sch_path: /headless/Documents/1bit_adc/3bit_dac.sch
**.subckt 3bit_dac ANALOG_IN SAR_SEL_0 SAR_SEL_1 SAR_SEL_2 IN1 OUT_DIGITAL NOUT_DIGITAL CLK RESET_B SET_B IN1
*.iopin ANALOG_IN
*.ipin SAR_SEL_0
*.ipin SAR_SEL_1
*.ipin SAR_SEL_2
*.iopin IN1
*.iopin OUT_DIGITAL
*.opin NOUT_DIGITAL
*.ipin CLK
*.ipin RESET_B
*.ipin SET_B
*.iopin IN1
XM1 ANALOG_IN SAR_SEL_0 net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VSS SAR_SEL_0 net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 ANALOG_IN SAR_SEL_1 net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 VSS SAR_SEL_1 net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 ANALOG_IN SAR_SEL_2 net3 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 VSS SAR_SEL_2 net3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR10 VR1 IN1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR1 net5 VR1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2 net2 net5 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR3 net6 VREF VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR4 net3 net6 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR5 net7 IN1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR6 net1 net7 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR7 VSS net8 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR8 VREF VR1 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
x1 net4 net4 IN1 net9 n_diffamp
XR9 VREF net9 VSS sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
**** begin user architecture code



.options gmin=1e-12
.option savecurrents
.option wnflag=1

.param vdd=1.8
.param clk=300n

VVDD VDD 0 DC {vdd}
VCLK CLK 0 PULSE(0 {vdd} 0 {clk/10} {clk/10} {1.5*clk} {2*clk})
VVSS VSS 0 DC 0
VVREF VREF 0 DC 3
VANALOG_IN 0 DC 0.9
VSET_B SET_B 0 DC {vdd}
VRESET_B RESET_B 0 DC {vdd}
*VSAR_SEL_2 SAR_SEL_2 0 0
*VSAR_SEL_1 SAR_SEL_1 0 0
*VSAR_SEL_0 SAR_SEL_0 0 0

*VANALOG_IN ANALOG_IN 0 pwl(0 0  0.5u 0.1  1u 0.2  1.5u 0.3  2u 0.4  2.5u 0.5  3u 0.6  3.5u 0.7  4u 0.8  4.5u 0.9  5u 1.0  5.5u 1.1  6u 1.2  6.5u 1.3  7u 1.4  7.5u 1.5  8u 1.6  8.5u 1.7  9u 1.8  9.5u 0  10u 0.1  10.5u 0.2  11u 0.3  11.5u 0.4  12u 0.5  12.5u 0.6  13u 0.7  13.5u 0.8  14u 0.9  14.5u 1.0  15u 1.1  15.5u 1.2  16u 1.3  16.5u 1.4  17u 1.5  17.5u 1.6  18u 1.7  18.5u 1.8  19u 0)
* Bit 0 (LSB) - period = 2us, toggles every 1us
VSAR_SEL_2 SAR_SEL_2 0 pwl(0 0  1u 0  1.1u 1.8  2u 1.8  2.1u 0  3u 0  3.1u 1.8  4u 1.8  4.1u 0  5u 0  5.1u 1.8  6u 1.8  6.1u 0  7u 0  7.1u 1.8  8u 1.8  8.1u 0  9u 0  9.1u 1.8  10u 1.8  10.1u 0  11u 0  11.1u 1.8  12u 1.8  12.1u 0  13u 0  13.1u 1.8  14u 1.8  14.1u 0  15u 0  15.1u 1.8  16u 1.8  16.1u 0  17u 0  17.1u 1.8  18u 1.8  18.1u 0  19u 0  19.1u 1.8  20u 1.8  20.1u 0  21u 0  21.1u 1.8  22u 1.8  22.1u 0  23u 0  23.1u 1.8  24u 1.8  24.1u 0  25u 0  25.1u 1.8  26u 1.8  26.1u 0  27u 0  27.1u 1.8  28u 1.8  28.1u 0  29u 0  29.1u 1.8  30u 1.8  30.1u 0  31u 0  31.1u 1.8  32u 1.8)
* Bit 1 - period = 4us, toggles every 2us
VSAR_SEL_1 SAR_SEL_1 0 pwl(0 0  2u 0  2.1u 1.8  4u 1.8  4.1u 0  6u 0  6.1u 1.8  8u 1.8  8.1u 0  10u 0  10.1u 1.8  12u 1.8  12.1u 0  14u 0  14.1u 1.8  16u 1.8  16.1u 0  18u 0  18.1u 1.8  20u 1.8  20.1u 0  22u 0  22.1u 1.8  24u 1.8  24.1u 0  26u 0  26.1u 1.8  28u 1.8  28.1u 0  30u 0  30.1u 1.8  32u 1.8)
* Bit 2 - period = 8us, toggles every 4us
VSAR_SEL_0 SAR_SEL_0 0 pwl(0 0  4u 0  4.1u 1.8  8u 1.8  8.1u 0  12u 0  12.1u 1.8  16u 1.8  16.1u 0  20u 0  20.1u 1.8  24u 1.8  24.1u 0  28u 0  28.1u 1.8  32u 1.8)
* Bit 3 (MSB) - period = 16us, toggles every 8us
VEN EN 0 pwl(0 0  8u 0  8.1u 1.8  16u 1.8  16.1u 0  24u 0  24.1u 1.8  32u 1.8)


.tran {clk/4} {clk*300}
.control

save all
echo TRAN
run
write 3bit_dac.raw all

.endc
.end



** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include /foss/pdks/sky130A/libs.tech/xschem/sky130_stdcells/

**** end user architecture code
**.ends

* expanding   symbol:  sky130_tests/n_diffamp.sym # of pins=4
** sym_path: /foss/pdks/volare/sky130/versions/0fe599b2afb6708d281543108caf8310912f54af/sky130A/libs.tech/xschem/sky130_tests/n_diffamp.sym
** sch_path: /foss/pdks/volare/sky130/versions/0fe599b2afb6708d281543108caf8310912f54af/sky130A/libs.tech/xschem/sky130_tests/n_diffamp.sch
.subckt n_diffamp OUT MINUS PLUS NBIAS
*.ipin PLUS
*.ipin MINUS
*.opin OUT
*.ipin NBIAS
XM1 net1 PLUS S GND sky130_fd_pr__nfet_01v8_lvt L=0.3 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT MINUS S GND sky130_fd_pr__nfet_01v8_lvt L=0.3 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.8 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.8 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 NBIAS GND GND sky130_fd_pr__nfet_01v8 L=1.2 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR1 GND S GND sky130_fd_pr__res_xhigh_po_0p35 L=50 mult=1 m=1
V5 S net2 0
.save i(v5)
.ends

.GLOBAL VSS
.GLOBAL VREF
.GLOBAL GND
.GLOBAL VDD
.end
