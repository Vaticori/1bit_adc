** sch_path: /headless/Documents/sar_adc/sar_adc/ideal_sar_adc.sch
**.subckt ideal_sar_adc
*  x3 -  sar_logic_analog  IS MISSING !!!!
vdd VDD GND 1.8
*  x1 -  ideal_comparator  IS MISSING !!!!
voffset net9 GND .6
vin net12 net9 sin(0 0.6 60 0)
C1 net10 GND 1p m=1
*  x2 -  ideal_dac  IS MISSING !!!!
*  x5 -  digital_to_real  IS MISSING !!!!
*  x6 -  ideal_ring_oscillator  IS MISSING !!!!
*  x7 -  ideal_bandgap_ref  IS MISSING !!!!
*  x4 -  transmission_gate  IS MISSING !!!!
v2 vin GND pulse(0 1.2 150us 25.6ms 0ns 100u 26ms)
**** begin user architecture code


.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.control
tran 100ns 30ms //16ms
plot v(digital_out_real) v(vin)
save all
run
write /foss/designs/sar_adc/ideal_sar_adc.raw
.endc




** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include /foss/pdks/sky130A/libs.tech/xschem/sky130_stdcells/
.include /headless/Documents/sar_adc/sar_adc/

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
