** sch_path: /headless/Documents/1bit_adc/passgate_2_outputs.sch
**.subckt passgate_2_outputs A OUT_1 OUT_0
*.ipin A
*.opin OUT_1
*.opin OUT_0
x1 OUT_1 net1 A net2 VDD VSS passgate W_N=1 L_N=0.2 W_P=1 L_P=0.2 m=1
x5 A VGND VNB VPB VPWR net2 sky130_fd_sc_hd__inv_1
x2 OUT_0 net3 net4 A VDD VSS passgate W_N=1 L_N=0.2 W_P=1 L_P=0.2 m=1
x3 A VGND VNB VPB VPWR net4 sky130_fd_sc_hd__inv_1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include /foss/pdks/sky130A/libs.tech/xschem/sky130_stdcells/

**** end user architecture code
**.ends

* expanding   symbol:  sky130_tests/passgate.sym # of pins=4
** sym_path: /foss/pdks/volare/sky130/versions/0fe599b2afb6708d281543108caf8310912f54af/sky130A/libs.tech/xschem/sky130_tests/passgate.sym
** sch_path: /foss/pdks/volare/sky130/versions/0fe599b2afb6708d281543108caf8310912f54af/sky130A/libs.tech/xschem/sky130_tests/passgate.sch
.subckt passgate Z A GP GN VCCBPIN VSSBPIN  W_N=1 L_N=0.2 W_P=1 L_P=0.2
*.iopin A
*.iopin Z
*.ipin GP
*.ipin GN
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
* noconn VCCBPIN
* noconn VSSBPIN
.ends

.end
